
module pll(
    input  wire osc_clk,
    output wire clk
    );

    assign clk = osc_clk;

endmodule
